`include "pipelined-mandelbrot";

module testbench ();
    
endmodule
